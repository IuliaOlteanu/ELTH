filtru trece-sus
vin 1 0 ac 1v pwl(0,0 0.2ms,0V 0.2001ms,1V 1ms, 1V)
R1 2 0 10
C1 1 2 15uF
.AC DEC 100 1Hz 100kHz
.tran 0.01ms 1ms
.probe
.end