Circuit cu STCC
R1 1 2 2
R2 2 4 1
R3 2 3 4
R5 5 0 2
V1 1 0 12
V3 5 3 4
I4 2 0 4
H2 4 5 V1 -2
.DC V1 12 12 1
.PRINT DC I(R1) I(R2) I(R3) I(R5) V(I4)
.END
