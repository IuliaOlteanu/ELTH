tema2
V1 3 5 50
V2 2 1 30
V3 0 5 90
R1 0 4 25
R2 2 5 12
R3 2 3 10
R4 0 1 10
R5 4 5 10
I1 3 4 2
.dc V3 90 90 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) I(V1) I(V2) I(V3) V(4,3) 
.end
