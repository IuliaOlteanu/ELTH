subpunctul c
R1 3 2 2
R2 4 0 2
R3 0 3 2
R4 0 1 2
V1 1 2 12
V2 3 4 6
G_curent 0 1 3 2 1
.DC V1 12 12 1
.PRINT DC I(R1) I(R2) I(R3) I(R4) V(G_curent)
.END
