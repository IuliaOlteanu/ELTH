tema1
V1 3 5 90
V2 0 5 50
V3 1 0 30
I1 3 4 6
R1 2 3 25
R2 4 5 12
R3 1 2 20
R4 2 5 10
R5 4 0 10
.dc V3 30 30 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) V(4,3) I(V2) I(V2) V(3) V(2) V(0) V(4) V(5)
.end
