Problema 1.3
V1 1 0 AC 40 45
V2 4 0 AC 80 45
R1 1 2 20
R2 2 5 10
L 5 0 31.841m
C 2 3 79.61u
R3 3 4 20
.AC LIN 1 50 50
.PRINT AC I(L) IP(L) I(R1) IP(R1) I(R2) IP(R2) I(R3) IP(R3) I(C) IP(C)
.END
