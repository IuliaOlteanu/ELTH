Problema 2
R1 1 2 610k
R2 3 0 10
R3 3 4 122000000
R4 5 0 15
L1 4 5 10m
C1 1 0 1/5u
V1 2 3 AC 14.14 -45
I1 5 2 AC 10 0
.AC LIN 1 0.159 0.159
.PRINT AC IR(V1) II(V1) IM(V1)
.END
