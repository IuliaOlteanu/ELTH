Problema 1.1
V1 1 0 AC 20 -45
L1 1 2 31.84M
L2 2 3 95.54M
R 3 4 10
V2 4 0 AC 60 45
C 2 0 159.15u
.AC LIN 1 50 50
.PRINT AC I(L1) IP(L1) I(R) IP(R) I(L2) IP(L2) I(C) IP(C)
.END
