Filtru trece-jos
Vin 1 0 AC 1
R 2 0 10k
C 1 2 10nF
.AC DEC 10 1hz 1meghz
.PROBE
.END
