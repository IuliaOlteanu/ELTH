regim tranzitoriu
c 0 3 100u ic=90
r2 3 0 10
l 3 0 62.5m ic=0
.tran 0.5ms 20ms uic
.probe
.end
