tema3
V1 0 4 90
V2 5 4 90
V3 2 4 50
R1 1 0 10
R2 2 1 5
R3 5 1 10
R4 0 3 30
R5 3 4 10
I1 2 3 5
.dc V1 90 90 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) I(V1) I(V2) I(V3) V(I1)
.end
