Aflarea conditiilor initiale
v1 2 1 90
r1 1 0 5
r2 3 0 10
c 2 3 100u
l 3 0 62.5m
.dc lin v1 90 90 1
.print dc v(2,3) i(l)
.end 

