simulare b)
V1 2 1 12
V2 2 3 24
R1 1 0 2
R2 3 4 8
R3 2 5 4
R4 4 5 4
R5 5 0 3
I1 0 4 3
.dc V1 12 12 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) V(I1)
.end
