fazori timp
V1 1 0 sin(0V 218.8V 50Hz 0 0 7.2)
V2 2 0 sin(0V 218.8V 50Hz 0 0 -112.8)
V3 3 0 sin(0V 218.8V 50Hz 0 0 127.2)
.tran 40ms 40ms 0 0.2ms
.probe
.end